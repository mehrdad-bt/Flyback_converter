** Profile: "Ideal_Devices-Tran"  [ D:\Work\Modelling\SMPS_DEsign_Kit\Demo_feb_12\AC_DC_VRM-PSpiceFiles\Ideal_Devices\Tran.sim ] 

** Creating circuit file "Tran.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../ac_dc_vrm-pspicefiles/ac_dc_vrm.lib" 
.LIB "../../../AC_DC_VRM-pspiceFiles/fwd_floating/tfrmr_subckt.lib" 
.LIB "../../../AC_DC_VRM-pspiceFiles/uc3843_test.lib" 
.LIB "../../../opto.lib" 
.LIB "../../../uc3843.lib" 
* From [PSPICE NETLIST] section of d:\Cadence\SPB_16.5\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 100m 0 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Ideal_Devices.net" 


.END
