** Profile: "Step_Load-step_current"  [ C:\ESD\Alok.Tri\cdssetup\OrCAD_Capture\16.6.0\tclscripts\caplearningresources\work\supportfiles\DesignExamples\SSFWDCNV\Designfiles\ssfwdcnv-pspicefiles\step_load\step_current.sim ] 

** Creating circuit file "step_current.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../ssfwdcnv-PSpiceFiles/ac_dc_vrm.lib" 
* From [PSPICE NETLIST] section of C:\ESD\Alok.Tri\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 20ms 10m 
.OPTIONS ADVCONV
.OPTIONS ABSTOL= 1.0n
.OPTIONS ITL4= 40
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) 
.INC "..\Step_Load.net" 


.END
